`timescale 1ns/1ps

module xnor_gate(input a, b, output y);
xnor(y, a, b);
endmodule
