`timescale 1ns/1ps

module buf_(input a, output y);
buf(y, a);
endmodule
