`timescale 1ns / 1ps

module or_gate(input a, b, output y);
or(y, a, b);
endmodule
