`timescale 1ns / 1ps
module not_gate(input a, output y);
not(y, a);
endmodule
